
module boot_code
(
    input  logic        CLK,
    input  logic        RSTN,

    input  logic        CSN,
    input  logic [9:0]  A,
    output logic [31:0] Q
  );

  const logic [0:547] [31:0] mem = {
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h00000013,
    32'h0100006F,
    32'h0100006F,
    32'h0080006F,
    32'h0040006F,
    32'h0000006F,
    32'h00000093,
    32'h00008113,
    32'h00008193,
    32'h00008213,
    32'h00008293,
    32'h00008313,
    32'h00008393,
    32'h00008413,
    32'h00008493,
    32'h00008513,
    32'h00008593,
    32'h00008613,
    32'h00008693,
    32'h00008713,
    32'h00008793,
    32'h00008813,
    32'h00008893,
    32'h00008913,
    32'h00008993,
    32'h00008A13,
    32'h00008A93,
    32'h00008B13,
    32'h00008B93,
    32'h00008C13,
    32'h00008C93,
    32'h00008D13,
    32'h00008D93,
    32'h00008E13,
    32'h00008E93,
    32'h00008F13,
    32'h00008F93,
    32'h00100117,
    32'hEF410113,
    32'h00001D17,
    32'h960D0D13,
    32'h00001D97,
    32'h958D8D93,
    32'h01BD5863,
    32'h000D2023,
    32'h004D0D13,
    32'hFFADDCE3,
    32'h00000513,
    32'h00000593,
    32'h076000EF,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h00000000,
    32'h46811101,
    32'h45A14601,
    32'h09F00513,
    32'h00EFCE06,
    32'h05134CE0,
    32'h00EF0400,
    32'h45815220,
    32'h00EF4501,
    32'h45815020,
    32'h00EF4501,
    32'h002854A0,
    32'h04000593,
    32'h58C000EF,
    32'h00812703,
    32'h01875513,
    32'h17B3157D,
    32'h0713DE87,
    32'h35332190,
    32'h886300A0,
    32'h670900E7,
    32'h8F990761,
    32'h00F037B3,
    32'h2083953E,
    32'h610501C1,
    32'h715D8082,
    32'hC6864505,
    32'hC2A6C4A2,
    32'hDE4EC0CA,
    32'hDA56DC52,
    32'hD65ED85A,
    32'hD266D462,
    32'h00EFD06A,
    32'h05933C20,
    32'h45010A10,
    32'h5AC000EF,
    32'h45014585,
    32'h2E0000EF,
    32'h45014585,
    32'h290000EF,
    32'h45014585,
    32'h338000EF,
    32'h87936785,
    32'hC0FBBB87,
    32'h00010037,
    32'h45810001,
    32'h00EF4501,
    32'h95373220,
    32'h45CD0000,
    32'h84450513,
    32'h5CC000EF,
    32'h27B74711,
    32'hC3D81A10,
    32'hF31FF0EF,
    32'h9537C911,
    32'h05930000,
    32'h05130250,
    32'h00EF8585,
    32'hA0015AE0,
    32'h00009537,
    32'h051345C9,
    32'h00EF8805,
    32'h45A159E0,
    32'h46014681,
    32'h00EF4519,
    32'h45013DE0,
    32'h434000EF,
    32'h45054581,
    32'h464000EF,
    32'h490000EF,
    32'h10055433,
    32'hFE143CE3,
    32'h80000637,
    32'h069345A1,
    32'h06130200,
    32'h05133486,
    32'h00EF0710,
    32'h45013AE0,
    32'h404000EF,
    32'h85224581,
    32'h434000EF,
    32'h460000EF,
    32'h10055533,
    32'hFE153CE3,
    32'h45214581,
    32'h3D0000EF,
    32'h02000693,
    32'h45A14601,
    32'h0EB00513,
    32'h37C000EF,
    32'h10000513,
    32'h3D0000EF,
    32'h45094581,
    32'h400000EF,
    32'h10000593,
    32'h00EF850A,
    32'h95374420,
    32'h45D90000,
    32'h89450513,
    32'h00C12C83,
    32'h2C034902,
    32'h24830041,
    32'h2A830101,
    32'h2B030141,
    32'h00EF01C1,
    32'h45814F20,
    32'h00EF4521,
    32'h5E6337A0,
    32'h64250790,
    32'h0C334981,
    32'h9BB7412C,
    32'h04130000,
    32'h9A378F04,
    32'h6D050000,
    32'h00891613,
    32'h02000693,
    32'h051345A1,
    32'h00EF0EB0,
    32'h652130A0,
    32'h360000EF,
    32'h45094581,
    32'h390000EF,
    32'h012C0533,
    32'h00EF65A1,
    32'h45993D20,
    32'h8ACB8513,
    32'h49C000EF,
    32'h0049D513,
    32'h95224585,
    32'h490000EF,
    32'hF649B533,
    32'h95224585,
    32'h484000EF,
    32'h45990985,
    32'h8B4A0513,
    32'h478000EF,
    32'h00EF996A,
    32'h91E34BE0,
    32'h00EFFB3C,
    32'h553337A0,
    32'h3CE31005,
    32'h9537FE15,
    32'h45B50000,
    32'h8BC50513,
    32'h454000EF,
    32'h49C000EF,
    32'h45214581,
    32'h2D8000EF,
    32'h07605E63,
    32'h89B36425,
    32'h4901409A,
    32'h00009BB7,
    32'h8F040413,
    32'h00009A37,
    32'h96136A85,
    32'h06930084,
    32'h45A10200,
    32'h0EB00513,
    32'h268000EF,
    32'h00EF6521,
    32'h45812BE0,
    32'h00EF4509,
    32'h85332EE0,
    32'h65A10099,
    32'h330000EF,
    32'h85134599,
    32'h00EF8ACB,
    32'h55133FA0,
    32'h45850049,
    32'h00EF9522,
    32'h35333EE0,
    32'h4585F649,
    32'h00EF9522,
    32'h09053E20,
    32'h05134599,
    32'h00EF8B4A,
    32'h94D63D60,
    32'h41C000EF,
    32'hFB2B11E3,
    32'h00009537,
    32'h02200593,
    32'h8CC50513,
    32'h3BC000EF,
    32'h404000EF,
    32'h1A1077B7,
    32'h0007A423,
    32'h08000793,
    32'h00078067,
    32'h00010001,
    32'h20830001,
    32'h450104C1,
    32'h04812403,
    32'h04412483,
    32'h04012903,
    32'h03C12983,
    32'h03812A03,
    32'h03412A83,
    32'h03012B03,
    32'h02C12B83,
    32'h02812C03,
    32'h02412C83,
    32'h02012D03,
    32'h80826161,
    32'h1A1076B7,
    32'h0006A783,
    32'hFF010113,
    32'h00F12623,
    32'h00100793,
    32'h00A797B3,
    32'h00C12703,
    32'hFFF7C793,
    32'h00E7F7B3,
    32'h00F12623,
    32'h00C12783,
    32'h00A595B3,
    32'h00F5E533,
    32'h00A12623,
    32'h00C12783,
    32'h00F6A023,
    32'h01010113,
    32'h00008067,
    32'h1A1017B7,
    32'h0007A783,
    32'hFF010113,
    32'h00F12623,
    32'h02058663,
    32'h00100713,
    32'h00C12783,
    32'h00A71533,
    32'h00F56533,
    32'h00A12623,
    32'h00C12703,
    32'h1A1017B7,
    32'h00E7A023,
    32'h01010113,
    32'h00008067,
    32'h00100793,
    32'h00A79533,
    32'hFFF54513,
    32'h00C12783,
    32'h00F57533,
    32'h00A12623,
    32'h00C12703,
    32'h1A1017B7,
    32'h00E7A023,
    32'h01010113,
    32'h00008067,
    32'h1A1017B7,
    32'hFF010113,
    32'h0087A783,
    32'h00F12623,
    32'h02058663,
    32'h00100713,
    32'h00C12783,
    32'h00A71533,
    32'h00F56533,
    32'h00A12623,
    32'h00C12703,
    32'h1A1017B7,
    32'h00E7A423,
    32'h01010113,
    32'h00008067,
    32'h00100793,
    32'h00A79533,
    32'hFFF54513,
    32'h00C12783,
    32'h00F57533,
    32'h00A12623,
    32'h00C12703,
    32'h1A1017B7,
    32'h00E7A423,
    32'h01010113,
    32'h00008067,
    32'hFF010113,
    32'h00812423,
    32'h00000593,
    32'h00050413,
    32'h00F00513,
    32'h00112623,
    32'hED1FF0EF,
    32'h00000593,
    32'h00E00513,
    32'hEC5FF0EF,
    32'h00000593,
    32'h00D00513,
    32'hEB9FF0EF,
    32'h00000593,
    32'h00C00513,
    32'hEADFF0EF,
    32'h04805663,
    32'h00000593,
    32'h01000513,
    32'hE9DFF0EF,
    32'h02142E63,
    32'h00000593,
    32'h00B00513,
    32'hE8DFF0EF,
    32'h02242663,
    32'h00000593,
    32'h00000513,
    32'hE7DFF0EF,
    32'h00342E63,
    32'h00C12083,
    32'h00812403,
    32'h00000593,
    32'h00100513,
    32'h01010113,
    32'hE61FF06F,
    32'h00C12083,
    32'h00812403,
    32'h01010113,
    32'h00008067,
    32'h00004837,
    32'hF0080813,
    32'h00869693,
    32'h02000713,
    32'h1A1027B7,
    32'h40B70733,
    32'h0106F6B3,
    32'hF265B5B3,
    32'h00E51533,
    32'h00878813,
    32'h00C78713,
    32'h00B6E5B3,
    32'h01078793,
    32'h00A82023,
    32'h00C72023,
    32'h00B7A023,
    32'h00008067,
    32'h01059593,
    32'h10055533,
    32'h00A5E5B3,
    32'h1A1027B7,
    32'h00B7AA23,
    32'h00008067,
    32'h1A102737,
    32'h01070713,
    32'h00072783,
    32'hFF010113,
    32'h00F12623,
    32'h00C12783,
    32'h1007D7B3,
    32'h01051513,
    32'h00F56533,
    32'h00A12623,
    32'h00C12783,
    32'h00F72023,
    32'h01010113,
    32'h00008067,
    32'h00100793,
    32'h00858593,
    32'h00B795B3,
    32'h00A79533,
    32'h000017B7,
    32'hF0078793,
    32'h00F5F5B3,
    32'hEE853533,
    32'h00A5E533,
    32'h1A1027B7,
    32'h00A7A023,
    32'h00008067,
    32'h1A1027B7,
    32'h0007A783,
    32'hFF010113,
    32'h00F12623,
    32'h00C12503,
    32'h01010113,
    32'h00008067,
    32'hD45597B3,
    32'hFF010113,
    32'hF455B5B3,
    32'h00F12423,
    32'h00058863,
    32'h00812783,
    32'h00178793,
    32'h00F12423,
    32'h00012623,
    32'h00C12683,
    32'h1A102737,
    32'h00812783,
    32'h02070813,
    32'h02F6DE63,
    32'h00072783,
    32'hCF0797B3,
    32'hFE078CE3,
    32'h00C12783,
    32'h00082583,
    32'h00C12683,
    32'h00168693,
    32'h00D12623,
    32'h01010613,
    32'h00279793,
    32'hFFC62603,
    32'h00812683,
    32'h00B567A3,
    32'hFCD646E3,
    32'h01010113,
    32'h00008067,
    32'h1A107737,
    32'h00470713,
    32'h00072603,
    32'h1A1007B7,
    32'hC0164633,
    32'h00C72023,
    32'h00478693,
    32'h00C78513,
    32'h0085D813,
    32'h08300713,
    32'h0FF5F593,
    32'h00E52023,
    32'h0106A023,
    32'h0A700713,
    32'h00B7A42B,
    32'h00E7A023,
    32'h00300793,
    32'h00F52023,
    32'h0006A783,
    32'h0F07F793,
    32'hC017C7B3,
    32'h00F6A023,
    32'h00008067,
    32'h04058263,
    32'h1A100637,
    32'h01460813,
    32'h00082783,
    32'h0207F793,
    32'hFE078CE3,
    32'h00150713,
    32'h0405468B,
    32'h1A1007B7,
    32'h00D7A023,
    32'hFFF58593,
    32'h03F450FB,
    32'h00058C63,
    32'h0017468B,
    32'hFFF58593,
    32'h00D62023,
    32'hFC0596E3,
    32'h00008067,
    32'h00008067,
    32'h1A100737,
    32'h01470713,
    32'h00072783,
    32'h0407F793,
    32'hFE078CE3,
    32'h00008067,
    32'h4C534953,
    32'h73274241,
    32'h6C757020,
    32'h6F6E6970,
    32'h000D0A21,
    32'h4F525245,
    32'h53203A52,
    32'h736E6170,
    32'h206E6F69,
    32'h20495053,
    32'h73616C66,
    32'h6F6E2068,
    32'h6F662074,
    32'h0A646E75,
    32'h0000000A,
    32'h64616F4C,
    32'h20676E69,
    32'h6D6F7266,
    32'h49505320};

  logic [9:0] A_Q;

  always_ff @(posedge CLK, negedge RSTN)
  begin
    if (~RSTN)
      A_Q <= '0;
    else
      if (~CSN)
        A_Q <= A;
  end

  assign Q = mem[A_Q];

endmodule